module rom_out(dout, addr);
	output [41:0] dout;
	input [7:0] addr;
	reg[41:0] mem[256:0];
	initial begin
	  /* mem[8'b00000000]=42'b1_00100_00000000_000_0_000000000000000001000011;	
		mem[8'b00000001]=42'b1_00100_00000001_000_0_000000000000000001000100;	//store
		//mem[8'b00000001]=42'b1_00001_00000000_000_0_000000000000000001000010;		//add
		mem[8'b00000010]=42'b1_00100_11111111_000_0_000000000000000000000000;	//store
	//	mem[8'b00000011]=42'b1_00001_00000000_000_0_000000000000000000000011; //add
		mem[8'b00000011]=42'b1_00011_11111111_000_0_000000000000000000000000;	//load
		mem[8'b00000100]=42'b0_00101_00000000_000_0_000000000000000000000000;  //outs
		mem[8'b00000101]=42'b1_00100_11111111_000_0_000000000000000000000001;	//store
		mem[8'b00000110]=42'b1_00011_11111111_000_0_000000000000000000000000;	//load
		mem[8'b00000111]=42'b0_00101_00000000_000_0_000000000000000000000000;  //outs
		*/
 		//$readmemb("/home/ryuji/Dropbox/elvm-cpu/rom.ecpu",mem);
		//$readmemb("C:/Users/ryuji/Dropbox/elvm-cpu/hello_rom.txt",mem);
		$readmemb("(place)/hello.ecpu",mem);

	end
	//rom memory(dout,addr,mem);
	assign dout = mem[addr];
endmodule
